program uvbot_main

   use shr_kind_mod,  only : r4 => shr_kind_r4

   use mpp_setup_mod,             only : mpp_init, mpp_end, mpp_barrier
   use mpp_setup_mod,             only : size, master, rank
   use mpp_io_mod,                only : error_handler, stdout
   use tprof_mod,                 only : tstart, tstop, tprnt

   use mpp_io_boundary_uvbot_mod, only : write_boundary_uvbot   
   use uvbot_mod,                 only : create_uvbot
   use uvbot_utils_mod,           only : uvbot_des_dims, uvbot_src_dims
   use uvbot_utils_mod,           only : uvbot_des_grid, uvbot_src_grid
   use time_mod,                  only : delt

   implicit none

   integer, parameter :: npx = 1
   integer, parameter :: npy = 1

   integer :: nxdes, nydes
   integer :: nxsrc, nysrc
   integer :: nrecs 

   real(KIND=r4), allocatable, dimension(:,:) :: uvbot_des
   real(KIND=r4), allocatable, dimension(:,:) :: uvbot_src

   real(KIND=r4), allocatable, dimension(:)   :: lon_des
   real(KIND=r4), allocatable, dimension(:)   :: lat_des

   real(KIND=r4), allocatable, dimension(:)   :: lon_src
   real(KIND=r4), allocatable, dimension(:)   :: lat_src

   real(KIND=r4) :: time_sec, time_hrs, time_day

   integer :: i, j, recs

   call mpp_init( npx, npy )

!  set size of destination grid
   call uvbot_des_dims ( nxdes, nydes )

!  set size of source grid  
   call uvbot_src_dims ( nxsrc, nysrc, nrecs )

!  allocate destination and source grids

   allocate ( uvbot_des(nxdes,nydes) )
   allocate ( uvbot_src(nxsrc,nysrc) )

   allocate ( lon_des(nxdes) )
   allocate ( lat_des(nydes) )

   allocate ( lon_src(nxsrc) )
   allocate ( lat_src(nysrc) )
  
!  set destination grid 
   call uvbot_des_grid ( uvbot_des, lon_des, lat_des, nxdes, nydes )

!  initialize uvbot_des fields

   call tstart('MAIN_UVBOT_LOOP')

   do recs=1,nrecs

     time_sec = (recs-1)*delt
     time_hrs = time_sec/3600.0
     time_day = time_hrs/24.0

!    set source grid 
     call uvbot_src_grid ( uvbot_src, lon_src, lat_src, nxsrc, nysrc, recs )

     write(stdout, 1000) recs
1000 format(2x, 'recs step = ', i4)

!    create interpolated fields

     call create_uvbot ( uvbot_src, uvbot_des, lon_src, lat_src, lon_des, lat_des, &
                                                        nxsrc, nysrc, nxdes, nydes )

     print *, MAXVAL(uvbot_des), MINVAL(uvbot_des)
     call write_boundary_uvbot ( uvbot_des, lon_des, lat_des, time_day, recs, &
                                                                 nxdes, nydes )

   enddo

   call tstop ('MAIN_UVBOT_LOOP')
   call tprnt

   call mpp_end

contains

end program uvbot_main

module mpp_io_boundary_model_spatial_mod

use shr_kind_mod,          only : r8 => shr_kind_r8
use shr_kind_mod,          only : r4 => shr_kind_r4
use mpp_setup_mod,         only : size, master, rank
use mpp_grid_mod,          only : mpp_get_global_indices
use mpp_io_mod,            only : get_unit_num, add_rank_to_file_name, error_handler
use mpp_io_mod,            only : stdout, read_diag_table
use mpp_update_domain_mod, only : update_domain

   implicit none
   private

   include 'netcdf.inc'

   public :: write_boundary_model_spatial

   logical :: first_time = .true.

   character(LEN=16), allocatable, dimension(:) :: diag_table_list
   integer :: num_diag_table

   character(LEN=48)  :: file_name ! file name associated with diags

   integer, parameter :: ndims_4d = 4 ! (i,j,k,t) dimensions in netCDF file
   integer, parameter :: ndims_3d = 3 ! (i,j,t)   dimensions in netCDF file

   integer :: start_4d(ndims_4d), count_4d(ndims_4d)
   integer :: start_3d(ndims_3d), count_3d(ndims_3d)

   character(LEN=32) :: var_units  ! units of variables

   character(LEN=32), parameter :: units   = 'units'
   character(LEN=32), parameter :: d_name  = 'domain_decomposition'

   character(LEN=32), parameter :: x_name    = 'x' ! name of x axis
   character(LEN=32), parameter :: y_name    = 'y' ! name of y axis
   character(LEN=32), parameter :: z_name    = 'z' ! name of z axis
   character(LEN=32), parameter :: rec_name  = 't' ! name of time axis

!  when we create netCDF files, variables and dimensions, we get back an ID for
!  each
   integer, dimension(ndims_4d) :: dimids_4d
   integer, dimension(ndims_3d) :: dimids_3d
   integer                      :: ncid, x_dimid, y_dimid, z_dimid, rec_dimid
   
   integer :: z_varid, y_varid, x_varid
 
   integer ::       um_varid,       vm_varid
   integer ::     ubot_varid,     vbot_varid
   integer ::     utop_varid,     vtop_varid
   integer ::     pgfx_varid,     pgfy_varid
   integer ::       wm_varid,      tur_varid
   integer ::     mask_varid,     znot_varid
   integer :: rain_acc_varid
  
contains
  
subroutine write_boundary_model_spatial ( um, vm, pgfx, pgfy, wm, tur, &
            znot, mask, rain_acc, recs, nx, ny, nz, ngx, ngy, npx, npy )

   integer, intent(in) :: nx, ny, nz
   integer, intent(in) :: ngx, ngy
   integer, intent(in) :: npx, npy

   real(KIND=r8) , dimension(:,:,:), intent(in)    :: um, vm
   real(KIND=r8) , dimension(:,:),   intent(inout) :: pgfx, pgfy
   real(KIND=r8) , dimension(:,:,:), intent(inout) :: wm, tur
   real(KIND=r8) , dimension(:,:),   intent(inout) :: znot, mask
   real(KIND=r8) , dimension(:,:),   intent(inout) :: rain_acc
   integer,                          intent(in)    :: recs
  
   real(kind=r8), dimension(ngx) :: xaxis
   real(kind=r8), dimension(ngy) :: yaxis
   real(kind=r8), dimension(nz)  :: zaxis
   
   real(KIND=r4), dimension(nx,ny,nz) :: var_write_4d_r4
   real(KIND=r4), dimension(nx,ny)    :: var_write_3d_r4

!  loop indexes, and error handling
   integer :: i, j, k, retval, id, io_unit

   integer :: mval(1)
   integer, parameter       :: nval = 4
   integer, dimension(nval) :: ival
   integer :: xbeg_data, xend_data, ybeg_data, yend_data
   integer :: xbeg_comp, xend_comp, ybeg_comp, yend_comp

   character(LEN=48) :: diag_file

   namelist /diagnostics/ diag_file

   if ( first_time == .true. ) then

!    set diags file names
     call get_unit_num (io_unit)
     open (io_unit,FILE='input.nml',STATUS='UNKNOWN')
     read (io_unit,NML=diagnostics)
     close(io_unit,STATUS='KEEP')

     if ( rank == master ) then
       write(stdout, 1000) diag_file
1000 format( 2x, 'name of diag file, written in: write_boundary_model_spatial = ', a48 )
     endif

     if ( npx*npy == 1 ) then
       file_name = diag_file
     else
       file_name = diag_file
       call add_rank_to_file_name(file_name)
     endif

!    read diag_table
     call read_diag_table ( diag_table_list, num_diag_table )

     id = rank + 1
     call mpp_get_global_indices ( xbeg_data, xend_data, ybeg_data, yend_data, &
                                   xbeg_comp, xend_comp, ybeg_comp, yend_comp, &
                                                id, nx, ny, ngx, ngy, npx, npy )

!    define axis 
     do k = 1, nz 
       zaxis(k) = k
     end do
     do j = 1, ngy
       yaxis(j) = j
     end do
     do i = 1, ngx
       xaxis(i) = i
     end do

!    create netCDF file, overwrite if already exists
     call write_boundary_model_state(1)

!    define the dimensions for each axis and get back ID for each
     retval = nf_def_dim(ncid, z_name  , nz                   , z_dimid  )
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_dim/z_dimid' )

     retval = nf_def_dim(ncid, y_name  , yend_data-ybeg_data+1, y_dimid  )
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_dim/y_dimid' )

     retval = nf_def_dim(ncid, x_name  , xend_data-xbeg_data+1, x_dimid  )
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_dim/x_dimid' )

     retval = nf_def_dim(ncid, rec_name, NF_UNLIMITED, rec_dimid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_dim/rec_dimid' )

!    define the coordinate variables
     retval = nf_def_var(ncid, z_name, NF_DOUBLE, 1, z_dimid, z_varid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/z_varid' )

     retval = nf_def_var(ncid, y_name, NF_DOUBLE, 1, y_dimid, y_varid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/y_varid' )

     retval = nf_def_var(ncid, x_name, NF_DOUBLE, 1, x_dimid, x_varid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/x_varid' )

     ival = (/1,ngx,xbeg_data,xend_data/)
     retval = NF_put_att_INT( ncid, x_varid, d_name, NF_INT, nval, ival )
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/NF_put_att_INT/ival' )

     ival = (/1,ngy,ybeg_data,yend_data/)
     retval = NF_put_att_INT( ncid, y_varid, d_name, NF_INT, nval, ival )
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/NF_put_att_INT/ival' )

     mval(1) = npx*npy
     retval = NF_PUT_ATT_INT( ncid, NF_GLOBAL, "NumFilesInSet", NF_INT, 1, mval ) 
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/NF_PUT_ATT_INT/mval' )

!    the dimids array is used to pass the ID of the dimensions of the
!    variables. Note that in fortran arrays are stored in column-major
     dimids_4d(1) = x_dimid
     dimids_4d(2) = y_dimid
     dimids_4d(3) = z_dimid
     dimids_4d(4) = rec_dimid

     dimids_3d(1) = x_dimid
     dimids_3d(2) = y_dimid
     dimids_3d(3) = rec_dimid

!    define the attributes for var
     do i=1,num_diag_table

       if ( TRIM(diag_table_list(i)) == 'ubot') then
         retval = nf_def_var(ncid, 'ubot'  , NF_REAL, ndims_3d, dimids_3d, ubot_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/ubot_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vbot') then
         retval = nf_def_var(ncid, 'vbot'  , NF_REAL, ndims_3d, dimids_3d, vbot_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/vbot_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'utop') then
         retval = nf_def_var(ncid, 'utop'  , NF_REAL, ndims_3d, dimids_3d, utop_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/utop_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vtop') then
         retval = nf_def_var(ncid, 'vtop'  , NF_REAL, ndims_3d, dimids_3d, vtop_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/vtop_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'um') then
         retval = nf_def_var(ncid, 'um'  , NF_REAL, ndims_4d, dimids_4d, um_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/um_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vm') then
         retval = nf_def_var(ncid, 'vm'  , NF_REAL, ndims_4d, dimids_4d, vm_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/vm_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'pgfx') then
         retval = nf_def_var(ncid, 'pgfx', NF_REAL, ndims_3d, dimids_3d, pgfx_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/pgfx_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'pgfy') then
         retval = nf_def_var(ncid, 'pgfy', NF_REAL, ndims_3d, dimids_3d, pgfy_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/pgfy_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'wm') then
         retval = nf_def_var(ncid, 'wm', NF_REAL, ndims_4d, dimids_4d, wm_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/wm_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'tur') then
         retval = nf_def_var(ncid, 'tur', NF_REAL, ndims_4d, dimids_4d, tur_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/tur_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'mask') then
         retval = nf_def_var(ncid, 'mask', NF_REAL, ndims_3d, dimids_3d, mask_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/mask_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'znot') then
         retval = nf_def_var(ncid, 'znot', NF_REAL, ndims_3d, dimids_3d, znot_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/znot_varid' )
       endif

       if ( TRIM(diag_table_list(i)) == 'rain_acc') then
         retval = nf_def_var(ncid, 'rain_acc', NF_REAL, ndims_3d, dimids_3d, rain_acc_varid)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_def_var/rain_acc_varid' )
       endif

       var_units = ''

       if ( TRIM(diag_table_list(i)) == 'ubot') then
         retval = nf_put_att_text(ncid, ubot_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vbot') then
         retval = nf_put_att_text(ncid, vbot_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'utop') then
         retval = nf_put_att_text(ncid, utop_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vtop') then
         retval = nf_put_att_text(ncid, vtop_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'um') then
         retval = nf_put_att_text(ncid, um_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'vm') then
         retval = nf_put_att_text(ncid, vm_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'pgfx') then
         retval = nf_put_att_text(ncid, pgfx_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif
  
       if ( TRIM(diag_table_list(i)) == 'pgfy') then
         retval = nf_put_att_text(ncid, pgfy_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif
 
       if ( TRIM(diag_table_list(i)) == 'wm') then
         retval = nf_put_att_text(ncid, wm_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'tur') then
         retval = nf_put_att_text(ncid, tur_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'mask') then
         retval = nf_put_att_text(ncid, mask_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif
  
       if ( TRIM(diag_table_list(i)) == 'znot') then
         retval = nf_put_att_text(ncid, znot_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

       if ( TRIM(diag_table_list(i)) == 'rain_acc') then
         retval = nf_put_att_text(ncid, rain_acc_varid, UNITS, len(var_units), var_units)
         if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_att_text/var_units' )
       endif

     enddo

!    end define mode; this tells netCDF we are done defining metadata
     retval = nf_enddef(ncid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_enddef' )

!    put axis data
     retval = nf_put_var_DOUBLE(ncid, z_varid, zaxis(1:nz))
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_DOUBLE/zaxis' )
  
     retval = nf_put_var_DOUBLE(ncid, y_varid, yaxis(ybeg_data:yend_data))
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_DOUBLE/yaxis' )
  
     retval = nf_put_var_DOUBLE(ncid, x_varid, xaxis(xbeg_data:xend_data))
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_DOUBLE/xaxis' )

     first_time = .false.
   else
!  open netCDF file
     call write_boundary_model_state(2)
   endif

   count_4d(1) = nx
   count_4d(2) = ny
   count_4d(3) = nz
   count_4d(4) = 1
   start_4d(1) = 1 
   start_4d(2) = 1 
   start_4d(3) = 1 
   start_4d(4) = recs

   count_3d(1) = nx
   count_3d(2) = ny
   count_3d(3) = 1
   start_3d(1) = 1 
   start_3d(2) = 1 
   start_3d(3) = recs

!  put var data 
   do i=1,num_diag_table

     if ( TRIM(diag_table_list(i)) == 'ubot') then
       var_write_3d_r4(:,:) = um(:,:,1)
       retval = nf_put_vara_REAL(ncid, ubot_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/ubot' )
     endif

     if ( TRIM(diag_table_list(i)) == 'vbot') then
       var_write_3d_r4(:,:) = vm(:,:,1)
       retval = nf_put_vara_REAL(ncid, vbot_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/vbot' )
     endif

     if ( TRIM(diag_table_list(i)) == 'utop') then
       var_write_3d_r4(:,:) = um(:,:,nz)
       retval = nf_put_vara_REAL(ncid, utop_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/utop' )
     endif

     if ( TRIM(diag_table_list(i)) == 'vtop') then
       var_write_3d_r4(:,:) = vm(:,:,nz)
       retval = nf_put_vara_REAL(ncid, vtop_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/vtop' )
     endif

     if ( TRIM(diag_table_list(i)) == 'um') then
       var_write_4d_r4(:,:,:) = um(:,:,:)
       retval = nf_put_vara_REAL(ncid, um_varid, start_4d, count_4d, var_write_4d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/um' )
     endif

     if ( TRIM(diag_table_list(i)) == 'vm') then
       var_write_4d_r4(:,:,:) = vm(:,:,:)
       retval = nf_put_vara_REAL(ncid, vm_varid, start_4d, count_4d, var_write_4d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/vm' )
     endif

     if ( TRIM(diag_table_list(i)) == 'pgfx') then
       call update_domain ( pgfx, nx, ny, npx, npy )
       var_write_3d_r4(:,:) = pgfx(:,:)
       retval = nf_put_vara_REAL(ncid, pgfx_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/pgfx' )
     endif

     if ( TRIM(diag_table_list(i)) == 'pgfy') then
       call update_domain ( pgfy, nx, ny, npx, npy )
       var_write_3d_r4(:,:) = pgfy(:,:)
       retval = nf_put_vara_REAL(ncid, pgfy_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/pgfy' )
     endif

     if ( TRIM(diag_table_list(i)) == 'wm') then
       var_write_4d_r4(:,:,:) = wm(:,:,:)
       retval = nf_put_vara_REAL(ncid, wm_varid, start_4d, count_4d, var_write_4d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/wm' )
     endif

     if ( TRIM(diag_table_list(i)) == 'tur') then
       var_write_4d_r4(:,:,:) = tur(:,:,:)
       retval = nf_put_vara_REAL(ncid, tur_varid, start_4d, count_4d, var_write_4d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/tur' )
     endif
     if ( TRIM(diag_table_list(i)) == 'mask') then
       call update_domain ( mask, nx, ny, npx, npy )
       var_write_3d_r4(:,:) = mask(:,:)
       retval = nf_put_vara_REAL(ncid, mask_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/mask' )
     endif

     if ( TRIM(diag_table_list(i)) == 'znot') then
       call update_domain ( znot, nx, ny, npx, npy )
       var_write_3d_r4(:,:) = znot(:,:)
       retval = nf_put_vara_REAL(ncid, znot_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/znot' )
     endif

     if ( TRIM(diag_table_list(i)) == 'rain_acc') then
       call update_domain ( rain_acc, nx, ny, npx, npy )
       var_write_3d_r4(:,:) = rain_acc(:,:)
       retval = nf_put_vara_REAL(ncid, rain_acc_varid, start_3d, count_3d, var_write_3d_r4)
       if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_spatial/nf_put_var_REAL/rain_acc' )
     endif

   enddo

   call write_boundary_model_state(3)

end subroutine write_boundary_model_spatial

subroutine write_boundary_model_state(case)
   integer, intent(in) :: case
   integer :: retval

   select CASE(case)
     CASE(1)
!    create netCDF file, overwrite if already exists
     retval = nf_create(file_name, nf_clobber, ncid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_state/nf_create' )

     CASE(2) 
!    open netCDF file
     retval = nf_open(file_name, nf_write, ncid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_state/nf_open' )

     CASE(3) 
!    close netCDF file
     retval = nf_close(ncid)
     if (retval .NE. 0) call error_handler ( 'ERROR', 'write_boundary_model_state/nf_close' )

    end select

end subroutine write_boundary_model_state

end module mpp_io_boundary_model_spatial_mod
